
module sign_ext(data_in, data_out);
	parameter WORD=8, EXT=4;
	input [WORD-1:0]data_in;
	output logic [WORD-1:0]data_out;
	
	
endmodule