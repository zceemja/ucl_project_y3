// Processor architecture
`define OISC
 
// Number of 16bit cells in ram 
`define RAM_SIZE 4096  

// Add debugging hardware to processor
`define DEBUG
