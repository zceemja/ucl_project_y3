// Processor architecture
`define OISC
 
// Number of 16bit cells in ram 
//`define RAM_SIZE 8192 
`define RAM_SIZE 4096

// Add debugging hardware to processor
`define DEBUG

`define ROMDIR "../../memory/build/"
`define RAMDIR "../../memory/build/"
